# LEF file generated for my_logo
VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO my_logo
   CLASS BLOCK ;
   FOREIGN my_logo 0 0 ;
   SIZE 120.000 BY 40.000 ;
   SYMMETRY X Y ;
   OBS
      LAYER met4 ;
         RECT 0.000 0.000 120.000 40.000 ;
      END
   END
END my_logo
