# LEF file generated for my_logo
VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

LAYER met4
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   PITCH 0.46 ;
   WIDTH 0.14 ;
   SPACING 0.14 ;
   RESISTANCE RPERSQ 0.0008 ;
   CAPACITANCE CPERSQDIST 0.00017 ;
   THICKNESS 0.14 ;
END met4

MACRO my_logo
   CLASS BLOCK ;
   FOREIGN my_logo 0 0 ;
   SIZE 80.000 BY 40.000 ;
   SYMMETRY X Y ;
   OBS
      LAYER met4 ;
         RECT 0.000 0.000 80.000 40.000 ;
      END
   END
END my_logo
